netcdf salinity_4 {
types:
  int(*) list_of_groups_t ;
  compound Metadata_t {
    int instrument ;
    byte manufacture ;
  }; // Metadata_t
dimensions:
	obs = 232323 ;
	copy = 3 ;
	qc_copy = 1 ;
variables:
	double time(obs) ;
		time:_FillValue = NaN ;
		time:long_name = "time of measurement" ;
		time:units = "seconds since 2001-07-01 12:33:24.000000" ;
		time:calendar = "gregorian" ;
	double lon(obs) ;
		lon:_FillValue = NaN ;
		lon:standard_name = "longitude" ;
		lon:long_name = "longitude of the observation" ;
		lon:units = "degrees_east" ;
	double lat(obs) ;
		lat:_FillValue = NaN ;
		lat:standard_name = "latitude" ;
		lat:long_name = "latitude of the observation" ;
		lat:units = "degrees_north" ;
	double vertical(obs) ;
		vertical:_FillValue = NaN ;
		vertical:long_name = "vertical distance above the surface" ;
		vertical:standard_name = "height" ;
		vertical:axis = "Z" ;
		vertical:ancillary_variables = "vertical_type" ;
	double observations(obs, copy) ;
		observations:_FillValue = NaN ;
		observations:long_name = "Observation data" ;
		observations:ancillary_variables = "error_variance truth obs_type" ;
		observations:coordinates = "lat lon vertical time" ;
	double error_variance(obs) ;
		error_variance:_FillValue = NaN ;
		error_variance:long_name = "error variance" ;
		error_variance:ancillary_variables = "obs_type" ;
		error_variance:coordinates = "lat lon vertical time" ;
	int qc(obs, qc_copy) ;
		qc:long_name = "quality control values" ;
		qc:ancillary_variables = "qc_copy" ;
		qc:flag_masks = 0, 1, 2, 3, 4, 5, 6 ;
		qc:flag_meanings = "assimilated evaluated assim_failed_postForwardOp eval_failed_postForwardOp unused_failed_priorForwardOp unselected failed_QC_check outlier" ;
		qc:coordinates = "lat lon vertical time" ;
	int qc_copy(qc_copy) ;
		qc_copy:long_name = "quality control types" ;
		qc_copy:flag_masks = 1, 2 ;
		qc_copy:flag_meanings = "Data_QC DART_QC" ;
	int obs_key(obs) ;
		obs_key:long_name = "DART key in linked list" ;
		obs_key:coordinates = "lat lon vertical time" ;
	list_of_groups_t list_of_groups(obs) ;
	Metadata_t Metadata(obs) ;
		Metadata:long_name = "Obseration Metadata" ;

// global attributes:
		:featureType = "point" ;
		:title = "Restructured netCDF file from Nancy" ;
		:author = "Jason Ngo, SIParCS Intern" ;
		:source = "Nancy Collins, NCAR|UCAR" ;
		:conventions = "CF-1.7" ;
		:creation_date = "YYYY MM DD HH MM SS = 2019 06 30 16 05 57" ;

group: Orange {
  variables:
  	int obs_id(obs) ;
  } // group Orange

group: Apple {
  variables:
  	int obs_id(obs) ;
  } // group Apple

group: Purple {
  variables:
  	int obs_id(obs) ;
  } // group Purple
}
