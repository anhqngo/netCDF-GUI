netcdf SOIL_SALINITY {
types:
//    int enum group_t {
//        Omega = 1, Oakton = 2, Plane = 3, Dummy = 4
//    };
    int(*) list_of_groups_t; // a variable-length array of group_id
//    compound Metadata_t {
//        int instrument;
//        list_of_groups_t list_of_groups;
//    }

dimensions:
    obs = 232323 ;
    copy = 3;
    qc_copy = 1;
variables:
	double time(obs) ;
		time:_FillValue = NaN ;
		time:long_name = "time of measurement" ;
		time:units = "seconds since 2001-07-01 12:33:24.000000" ;
		time:calendar = "gregorian" ;
	double lon(obs) ;
		lon:_FillValue = NaN ;
		lon:standard_name = "longitude" ;
		lon:long_name = "longitude of the observation" ;
		lon:units = "degrees_east" ;
	double lat(obs) ;
		lat:_FillValue = NaN ;
		lat:standard_name = "latitude" ;
		lat:long_name = "latitude of the observation" ;
		lat:units = "degrees_north" ;
	double vertical(obs) ;
		vertical:_FillValue = NaN ;
		vertical:long_name = "vertical distance above the surface" ;
		vertical:standard_name = "height" ;
		vertical:axis = "Z" ;

	double observation(obs,copy) ;
		observation:_FillValue = NaN ;
		observation:long_name = "Observation data" ;
		observation:ancillary_variables = "Metadata" ;
		observation:coordinates = "lat lon vertical time" ;

	int qc(obs, qc_copy) ;
		qc:long_name = "quality control values" ;
		qc:ancillary_variables = "qc_copy" ;
		qc:flag_masks = 0, 1, 2, 3, 4, 5, 6 ;
		qc:flag_meanings = "assimilated evaluated assim_failed_postForwardOp eval_failed_postForwardOp unused_failed_priorForwardOp unselected failed_QC_check outlier" ;
		qc:coordinates = "lat lon vertical time" ;
	int qc_copy(qc_copy) ;
		qc_copy:long_name = "quality control types" ;
		qc_copy:flag_masks = 1, 2 ;
		qc_copy:flag_meanings = "Data_QC DART_QC" ;

    list_of_groups_t list_of_groups(obs);

//    Metadata_t Metadata(obs);

// global attributes:
		:featureType = "point" ;
		:title = "Restructured netCDF file from Tim" ;
		:author = "Jason Ngo, SIParCS Intern" ;
		:source = "Tim Hoar, NCAR|UCAR" ;
		:conventions = "CF-1.7" ;
		:creation_date = "YYYY MM DD HH MM SS = 2019 07 08 16 05 57" ;

data:
    time = 500, 600;
    lat = 50, 80;
    lon = 30, 80;
    vertical = 3, 3;
    list_of_groups = {1}, {1,2};
//    Metadata = {_, _}, {_,_};

//  groups:
    group: Europe {
        variables:
            int obs_id(obs);
        data: 
            obs_id = 1; // Pointer to the observation data
    }
    group: Apple_manufacture {
        variables:
            int obs_id(obs);
        data: 
            obs_id = 1, 2; // Pointer to the observation data
    }
}
